library ieee;
use ieee.std_logic_1164.all;
use work.testing_functions.all;
use work.data_link_pkg.all;

entity ilas_parser_tb is
end entity ilas_parser_tb;

architecture a1 of ilas_parser_tb is
  type test_vector is record
    ci_state : link_state;
    di_char  : link_character;

    expected_finished : std_logic;
    expected_error : std_logic;
    expected_wrong_chksum : std_logic;
    expected_unexpected_char : std_logic;
    expected_config_index : integer;
  end record test_vector;

  type config_array is array (natural range<>) of link_config;
  constant config_vectors : config_array :=
  (
    (
      DID => 170,
      ADJCNT =>  7,
      BID => 14,
      ADJDIR => '1',
      PHADJ => '1',
      LID => 10,
      SCR => '1',
      L => 31,
      F => 205,
      K => 32,
      M => 52,
      CS => 2,
      N => 4,
      SUBCLASSV => 1,
      Nn => 30,
      JESDV => 0,
      S => 1,
      HD => '0',
      CF =>  0,
      RES1 => "11111111",
      RES2 => "00000000",
      X => "010010000",
      CHKSUM => 48
    ),
    (
      DID => 170,
      ADJCNT =>  7,
      BID => 14,
      ADJDIR => '1',
      PHADJ => '1',
      LID => 10,
      SCR => '1',
      L => 31,
      F => 205,
      K => 32,
      M => 52,
      CS => 2,
      N => 4,
      SUBCLASSV => 1,
      Nn => 30,
      JESDV => 0,
      S => 1,
      HD => '0',
      CF =>  0,
      RES1 => "11111111",
      RES2 => "11111111",
      X => "010010000",
      CHKSUM => 48
    )
  );

  type test_vector_array is array (natural range<>) of test_vector;
  constant test_vectors : test_vector_array :=
  (
    -- correct sequence, config index 0
    (INIT, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (CGS,  ('1', '0', '0', "10111100", '0'), '0', '0', '0', '0', -1),
    (CGS,  ('1', '0', '0', "10111100", '0'), '0', '0', '0', '0', -1),
    (CGS,  ('1', '0', '0', "10111100", '0'), '0', '0', '0', '0', -1),
    (CGS,  ('1', '0', '0', "10111100", '0'), '0', '0', '0', '0', -1),
    (ILS, ('1', '0', '0', "00011100", '0'), '0', '0', '0', '0', -1),  -- R, 0 mult
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('1', '0', '0', "01111100", '0'), '0', '0', '0', '0', -1),  -- A
    (ILS, ('1', '0', '0', "00011100", '0'), '0', '0', '0', '0', -1),  -- R, 1 mult
    (ILS, ('1', '0', '0', "10011100", '0'), '0', '0', '0', '0', -1),  -- 28.4
    (ILS, ('0', '0', '0', "10101010", '0'), '0', '0', '0', '0', -1),  -- DID
    (ILS, ('0', '0', '0', "01111110", '0'), '0', '0', '0', '0', -1),  -- ADJCNT,BID
    (ILS, ('0', '0', '0', "01101010", '0'), '0', '0', '0', '0', -1),  -- X,ADJDIR,PHADJ,LID
    (ILS, ('0', '0', '0', "11011110", '0'), '0', '0', '0', '0', -1),  -- SCR,X,L
    (ILS, ('0', '0', '0', "11001100", '0'), '0', '0', '0', '0', -1),  -- F
    (ILS, ('0', '0', '0', "01011111", '0'), '0', '0', '0', '0', -1),  -- X, K
    (ILS, ('0', '0', '0', "00110011", '0'), '0', '0', '0', '0', -1),  -- M
    (ILS, ('0', '0', '0', "10000011", '0'), '0', '0', '0', '0', -1),  -- CS,X,N
    (ILS, ('0', '0', '0', "00111101", '0'), '0', '0', '0', '0', -1),  -- SUBCLASSV,Nn
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),  -- JESDV,S
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "11111111", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00110000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('1', '0', '0', "01111100", '0'), '0', '0', '0', '0',  0),  -- A
    (ILS, ('1', '0', '0', "00011100", '0'), '0', '0', '0', '0',  0),  -- R
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('1', '0', '0', "01111100", '0'), '0', '0', '0', '0',  0),  -- A
    (ILS, ('1', '0', '0', "00011100", '0'), '0', '0', '0', '0',  0),  -- R, 2 mult
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0',  0),
    (ILS, ('1', '0', '0', "01111100", '0'), '1', '0', '0', '0',  0),  -- A
    (DATA, ('0', '0', '0', "00000001", '0'), '1', '0', '0', '0',  0),
    (DATA, ('0', '0', '0', "00000010", '0'), '1', '0', '0', '0',  0),
    (DATA, ('0', '0', '0', "00000011", '0'), '1', '0', '0', '0',  0),
    -- incorrect sequence - /R/ at wrong place
    (INIT, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (CGS,  ('1', '0', '0', "10111100", '0'), '0', '0', '0', '0', -1),
    (CGS,  ('1', '0', '0', "10111100", '0'), '0', '0', '0', '0', -1),
    (CGS,  ('1', '0', '0', "10111100", '0'), '0', '0', '0', '0', -1),
    (CGS,  ('1', '0', '0', "10111100", '0'), '0', '0', '0', '0', -1),
    (ILS, ('1', '0', '0', "00011100", '0'), '0', '0', '0', '0', -1),  -- R, 0 mult
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('1', '0', '0', "00011100", '0'), '0', '1', '0', '1', -1),  -- R, wrong place
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '1', '0', '1', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '1', '0', '1', -1),
    (INIT, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    -- incorrect sequence - /A/ at wrong place
    (INIT, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (CGS,  ('1', '0', '0', "10111100", '0'), '0', '0', '0', '0', -1),
    (CGS,  ('1', '0', '0', "10111100", '0'), '0', '0', '0', '0', -1),
    (CGS,  ('1', '0', '0', "10111100", '0'), '0', '0', '0', '0', -1),
    (CGS,  ('1', '0', '0', "10111100", '0'), '0', '0', '0', '0', -1),
    (ILS, ('1', '0', '0', "00011100", '0'), '0', '0', '0', '0', -1),  -- R, 0 mult
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('1', '0', '0', "01111100", '0'), '0', '1', '0', '1', -1),  -- A
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '1', '0', '1', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '1', '0', '1', -1),
    (INIT, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    -- incorrect sequence - wrong check sum
    (INIT, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (CGS,  ('1', '0', '0', "10111100", '0'), '0', '0', '0', '0', -1),
    (CGS,  ('1', '0', '0', "10111100", '0'), '0', '0', '0', '0', -1),
    (CGS,  ('1', '0', '0', "10111100", '0'), '0', '0', '0', '0', -1),
    (CGS,  ('1', '0', '0', "10111100", '0'), '0', '0', '0', '0', -1),
    (ILS, ('1', '0', '0', "00011100", '0'), '0', '0', '0', '0', -1),  -- R, 0 mult
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('1', '0', '0', "01111100", '0'), '0', '0', '0', '0', -1),  -- A
    (ILS, ('1', '0', '0', "00011100", '0'), '0', '0', '0', '0', -1),  -- R, 1 mult
    (ILS, ('1', '0', '0', "10011100", '0'), '0', '0', '0', '0', -1),  -- 28.4
    (ILS, ('0', '0', '0', "10101010", '0'), '0', '0', '0', '0', -1),  -- DID
    (ILS, ('0', '0', '0', "01111110", '0'), '0', '0', '0', '0', -1),  -- ADJCNT,BID
    (ILS, ('0', '0', '0', "01001010", '0'), '0', '0', '0', '0', -1),  -- X,ADJDIR,PHADJ,LID
    (ILS, ('0', '0', '0', "11011110", '0'), '0', '0', '0', '0', -1),  -- SCR,X,L
    (ILS, ('0', '0', '0', "11001100", '0'), '0', '0', '0', '0', -1),  -- F
    (ILS, ('0', '0', '0', "01011111", '0'), '0', '0', '0', '0', -1),  -- X, K
    (ILS, ('0', '0', '0', "00110011", '0'), '0', '0', '0', '0', -1),  -- M
    (ILS, ('0', '0', '0', "10000011", '0'), '0', '0', '0', '0', -1),  -- CS,X,N
    (ILS, ('0', '0', '0', "00111101", '0'), '0', '0', '0', '0', -1),  -- SUBCLASSV,Nn
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),  -- JESDV,S
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "11111111", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '0', '0', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '1', '1', '0', -1),
    (ILS, ('1', '0', '0', "01111100", '0'), '0', '1', '1', '0', -1),  -- A
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '1', '1', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '1', '1', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '1', '1', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '1', '1', '0', -1),
    (ILS, ('0', '0', '0', "00000000", '0'), '0', '1', '1', '0', -1),
    (INIT, ('0', '0', '0', "00000000", '0'), '0', '1', '1', '0', -1)
  );

  constant clk_period : time := 1 ns;

  constant F : integer range 0 to 256 := 17;
  constant K : integer range 0 to 32 := 1;

  signal clk : std_logic := '0';
  signal reset : std_logic := '0';

  signal ci_state : link_state := INIT;

  signal di_char : link_character;
  signal do_config : link_config;

  signal co_finished : std_logic;
  signal co_error : std_logic;
  signal co_wrong_chksum : std_logic;
  signal co_unexpected_char : std_logic;

  signal test_data_index : integer := 0;

begin  -- architecture a1
  uut: entity work.ilas_parser
    generic map (
      F => F,
      K => K)
    port map (
      ci_char_clk => clk,
      ci_reset    => reset,
      ci_state    =>  ci_state,
      di_char     => di_char,
      do_config   => do_config,
      co_finished => co_finished,
      co_error    => co_error,
      co_wrong_chksum    => co_wrong_chksum,
      co_unexpected_char => co_unexpected_char);

  clk_gen: process is
  begin -- process clk_gen
    wait for clk_period/2;
	 clk <= not clk;
  end process clk_gen;
  
  reset_gen: process is
  begin -- process reset_gen
    wait for clk_period*2;
    reset <= '1';
  end process reset_gen;

  test: process is
    variable test_vec : test_vector;
    variable prev_test_vec : test_vector;
  begin  -- process test
    wait for clk_period*2;

    for i in test_vectors'range loop
      test_data_index <= i;
      test_vec := test_vectors(i);
      di_char <= test_vec.di_char;
      ci_state <= test_vec.ci_state;

      if i > 0 then
        prev_test_vec := test_vectors(i - 1);

        if prev_test_vec.expected_config_index > -1 then
        assert do_config = config_vectors(prev_test_vec.expected_config_index) report "The config does not match. Index: " & integer'image(i-1) severity error;
        end if;

        assert co_error = prev_test_vec.expected_error report "The error does not match. Index: " & integer'image(i-1) severity error;
        assert co_wrong_chksum = prev_test_vec.expected_wrong_chksum report "The wrong_chksum does not match. Index: " & integer'image(i-1) severity error;
        assert co_unexpected_char = prev_test_vec.expected_unexpected_char report "The unexpected_char does not match. Index: " & integer'image(i-1) severity error;
        assert co_finished = prev_test_vec.expected_finished report "The finished does not match. Index: " & integer'image(i-1) severity error;
      end if;

      wait for clk_period;
    end loop;  -- i
    wait for 100 ms;
  end process test;
end architecture a1;
