library ieee;
use ieee.std_logic_1164.all;
use work.testing_functions.all;
use work.data_link_pkg.all;

entity ilas_parser_tb is
end entity ilas_parser_tb;

architecture a1 of ilas_parser_tb is
  type test_vector is record
    ci_state : link_state;
    di_char  : character_vector;

    expected_finished : std_logic;
    expected_error : std_logic;
    expected_wrong_chksum : std_logic;
    expected_unexpected_char : std_logic;
    expected_config_index : integer;
  end record test_vector;

  type config_array is array (natural range<>) of link_config;
  constant config_vectors : config_array :=
  (
    -- DID = 10101010
    -- ADJCNT = 0111
    -- BID = 1110
    -- ADJDIR = 1
    -- PHADJ = 0
    -- LID 01010
    -- SCR = 1
    -- L = 11110
    -- F = 11001100
    -- K = 11111
    -- M = 00110011
    -- CS = 10
    -- N = 00011
    -- SUBCLASSV = 1
    -- Nn = 11101
    -- JESDV = 0
    -- S = 0
    -- HD = 0
    -- CF = 0
    -- RES1 = 11111111
    -- RES2 = 00000000
    -- X = 010010000
  );

  type test_vector_array is array (natural range<>) of test_vector;
  constant test_vectors : test_vector_array :=
  (
    -- correct sequence, config index 0
    (INIT, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (CGS,  ('0', '0', '0', "10111100"), '0', '0', '0', '0', -1),
    (CGS,  ('0', '0', '0', "10111100"), '0', '0', '0', '0', -1),
    (CGS,  ('0', '0', '0', "10111100"), '0', '0', '0', '0', -1),
    (CGS,  ('0', '0', '0', "10111100"), '0', '0', '0', '0', -1),
    (ILAS, ('1', '0', '0', "00011100"), '0', '0', '0', '0', -1),  -- R, 0 mult
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('1', '0', '0', "01111100"), '0', '0', '0', '0', -1),  -- A
    (ILAS, ('1', '0', '0', "00011100"), '0', '0', '0', '0', -1),  -- R, 1 mult
    (ILAS, ('1', '0', '0', "10011100"), '0', '0', '0', '0', -1),  -- 28.4
    (ILAS, ('0', '0', '0', "10101010"), '0', '0', '0', '0', -1),  -- DID
    (ILAS, ('0', '0', '0', "01111110"), '0', '0', '0', '0', -1),  -- ADJCNT,BID
    (ILAS, ('0', '0', '0', "01001010"), '0', '0', '0', '0', -1),  -- X,ADJDIR,PHADJ,LID
    (ILAS, ('0', '0', '0', "11011110"), '0', '0', '0', '0', -1),  -- SCR,X,L
    (ILAS, ('0', '0', '0', "11001100"), '0', '0', '0', '0', -1),  -- F
    (ILAS, ('0', '0', '0', "01011111"), '0', '0', '0', '0', -1),  -- X, K
    (ILAS, ('0', '0', '0', "00110011"), '0', '0', '0', '0', -1),  -- M
    (ILAS, ('0', '0', '0', "10000011"), '0', '0', '0', '0', -1),  -- CS,X,N
    (ILAS, ('0', '0', '0', "00111101"), '0', '0', '0', '0', -1),  -- SUBCLASSV,Nn
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),  -- JESDV,S
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "11111111"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00110000"), '0', '0', '0', '0', -1),
    (ILAS, ('1', '0', '0', "01111100"), '0', '0', '0', '0',  0),  -- A
    (ILAS, ('1', '0', '0', "00011100"), '0', '0', '0', '0',  0),  -- R
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('1', '0', '0', "01111100"), '0', '0', '0', '0',  0),  -- A
    (ILAS, ('1', '0', '0', "00011100"), '0', '0', '0', '0',  0),  -- R, 2 mult
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0',  0),
    (ILAS, ('1', '0', '0', "01111100"), '0', '0', '0', '0',  0),  -- A
    (DATA, ('0', '0', '0', "00000001"), '1', '0', '0', '0',  0),
    (DATA, ('0', '0', '0', "00000010"), '1', '0', '0', '0',  0),
    (DATA, ('0', '0', '0', "00000011"), '1', '0', '0', '0',  0),
    -- incorrect sequence - /R/ at wrong place
    (INIT, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (CGS,  ('0', '0', '0', "10111100"), '0', '0', '0', '0', -1),
    (CGS,  ('0', '0', '0', "10111100"), '0', '0', '0', '0', -1),
    (CGS,  ('0', '0', '0', "10111100"), '0', '0', '0', '0', -1),
    (CGS,  ('0', '0', '0', "10111100"), '0', '0', '0', '0', -1),
    (ILAS, ('1', '0', '0', "00011100"), '0', '0', '0', '0', -1),  -- R, 0 mult
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('1', '0', '0', "00011100"), '0', '1', '0', '1', -1),  -- R, wrong place
    (ILAS, ('0', '0', '0', "00000000"), '0', '1', '0', '1', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '1', '0', '1', -1),
    (INIT, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    -- incorrect sequence - /A/ at wrong place
    (INIT, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (CGS,  ('0', '0', '0', "10111100"), '0', '0', '0', '0', -1),
    (CGS,  ('0', '0', '0', "10111100"), '0', '0', '0', '0', -1),
    (CGS,  ('0', '0', '0', "10111100"), '0', '0', '0', '0', -1),
    (CGS,  ('0', '0', '0', "10111100"), '0', '0', '0', '0', -1),
    (ILAS, ('1', '0', '0', "00011100"), '0', '0', '0', '0', -1),  -- R, 0 mult
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('1', '0', '0', "01111100"), '0', '1', '0', '1',  0),  -- A
    (ILAS, ('0', '0', '0', "00000000"), '0', '1', '0', '1', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '1', '0', '1', -1),
    (INIT, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    -- incorrect sequence - wrong check sum
    (INIT, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (CGS,  ('0', '0', '0', "10111100"), '0', '0', '0', '0', -1),
    (CGS,  ('0', '0', '0', "10111100"), '0', '0', '0', '0', -1),
    (CGS,  ('0', '0', '0', "10111100"), '0', '0', '0', '0', -1),
    (CGS,  ('0', '0', '0', "10111100"), '0', '0', '0', '0', -1),
    (ILAS, ('1', '0', '0', "00011100"), '0', '0', '0', '0', -1),  -- R, 0 mult
    (ILAS, ('1', '0', '0', "00011100"), '0', '0', '0', '0', -1),  -- R, 0 mult
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('1', '0', '0', "01111100"), '0', '0', '0', '0', -1),  -- A
    (ILAS, ('1', '0', '0', "00011100"), '0', '0', '0', '0', -1),  -- R, 1 mult
    (ILAS, ('1', '0', '0', "10011100"), '0', '0', '0', '0', -1),  -- 28.4
    (ILAS, ('0', '0', '0', "10101010"), '0', '0', '0', '0', -1),  -- DID
    (ILAS, ('0', '0', '0', "01111110"), '0', '0', '0', '0', -1),  -- ADJCNT,BID
    (ILAS, ('0', '0', '0', "01001010"), '0', '0', '0', '0', -1),  -- X,ADJDIR,PHADJ,LID
    (ILAS, ('0', '0', '0', "11011110"), '0', '0', '0', '0', -1),  -- SCR,X,L
    (ILAS, ('0', '0', '0', "11001100"), '0', '0', '0', '0', -1),  -- F
    (ILAS, ('0', '0', '0', "01011111"), '0', '0', '0', '0', -1),  -- X, K
    (ILAS, ('0', '0', '0', "00110011"), '0', '0', '0', '0', -1),  -- M
    (ILAS, ('0', '0', '0', "10000011"), '0', '0', '0', '0', -1),  -- CS,X,N
    (ILAS, ('0', '0', '0', "00111101"), '0', '0', '0', '0', -1),  -- SUBCLASSV,Nn
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),  -- JESDV,S
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "11111111"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '0', '0', '0', -1),
    (ILAS, ('1', '0', '0', "01111100"), '0', '1', '1', '0', -1),  -- A
    (ILAS, ('0', '0', '0', "00000000"), '0', '1', '1', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '1', '1', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '1', '1', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '1', '1', '0', -1),
    (ILAS, ('0', '0', '0', "00000000"), '0', '1', '1', '0', -1)
  );

  constant clk_period : time := 1 ns;

  constant F : integer range 0 to 256 := 17;

  signal clk : std_logic := '0';
  signal reset : std_logic := '0';

  signal ci_state : link_state := INIT;

  signal di_char : character_vector;
  signal do_config : link_config;

  signal co_finished : std_logic;
  signal co_error : std_logic;
  signal co_wrong_chksum : std_logic;
  signal co_unexpected_char : std_logic;

  signal test_data_index : integer := 0;

begin  -- architecture a1
  uut: entity work.ilas_parser
    port map (
      ci_char_clk => clk,
      ci_reset    => reset,
      ci_F        => F,
      ci_state    =>  ci_state,
      di_char     => di_char,
      do_config   => do_config,
      co_finished => co_finished,
      co_error    => co_error,
      co_wrong_chksum    => co_wrong_chksum,
      co_unexpected_char => co_unexpected_char);

  clk <= not clk after clk_period/2;
  reset <= '1' after clk_period*2;

  test: process is
    variable test_vec : test_vector;
    variable prev_test_vec : test_vector;
  begin  -- process test
    wait for clk_period*2;

    for i in test_vectors'range loop
      test_data_index <= i;
      test_vec := test_vectors(i);
      di_char <= test_vec.di_char;
      ci_state <= test_vec.ci_state;

      if i > 0 then
        prev_test_vec := test_vectors(i - 1);

        if prev_test_vec.expected_config_index > -1 then
          assert co_config = config_vectors(prev_test_vec.expected_config_index) report "The config does not match. Index: " & integer'image(i-1) severity error;
        end if;

        assert co_error = prev_test_vec.expected_error report "The error does not match. Index: " & integer'image(i-1) severity error;
        assert co_wrong_chksum = prev_test_vec.expected_wrong_chksum report "The wrong_chksum does not match. Index: " & integer'image(i-1) severity error;
        assert co_unexpected_char = prev_test_vec.expected_unexpected_char report "The unexpected_char does not match. Index: " & integer'image(i-1) severity error;
        assert co_finished = prev_test_vec.expected_finished report "The finished does not match. Index: " & integer'image(i-1) severity error;
      end if;

      wait for clk_period;
    end loop;  -- i
    wait for 100 ms;
  end process test;
end architecture a1;
